module dddd (
    input clk
);
    
endmodule