module dddd (
    input clk,
    input rst
);
    
endmodule