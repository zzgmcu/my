module dddd (
    input clk,
    input rst,
    output c
);
    
endmodule